ENTITY app IS
END ENTITY;

ARCHITECTURE rtl OF app IS
BEGIN
END ARCHITECTURE;